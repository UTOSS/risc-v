`ifndef PARAMS_VH
`define PARAMS_VH

//Opcodes
parameter RType = 7'b0110011
parameter IType = 7'b0010011 //excluding lw 
parameter LWType = 7'b0000011
parameter SType = 7'b0100011
parameter BType = 7'b1100011
parameter JType = 7'b1101111

`endif // PARAMS_VH
