`ifndef PARAMS_VH
`define PARAMS_VH

`endif // PARAMS_VH