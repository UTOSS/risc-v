`timescale 1ns/1ps

`include "src/types.svh"      // <-- bring in enum literals like PC_SRC__JUMP
`include "test/utils.svh"

/* verilator lint_off IMPORTSTAR */
/* verilator lint_off UNUSEDSIGNAL */
/* verilator lint_off INITIALDLY */

import pkg_control_fsm::*;

module jal_tb;

  reg clk;
  reg reset;

  // DUT
  top uut
    ( .clk   ( clk   )
    , .reset ( reset )
    );

  // 10ns clock
  initial begin
    clk = 0;
    forever #5 clk = ~clk;
  end

  // helper: wait one cycle then assert expected FSM state
  /* verilator lint_off UNUSEDSIGNAL */
  task wait_till_next_cfsm_state(input state_t expected_state);
  /* verilator lint_on UNUSEDSIGNAL */
    @(posedge clk); #1;
    `assert_equal(uut.core.control_fsm.current_state, expected_state)
  endtask

  initial begin
    reset = `TRUE;

    // Program:
    //   0x00000000: JAL x1, +16   (target = 16)
    // J-type encoding: opcode=0x6F, rd=x1, imm=+16 -> 0x010000EF
    uut.memory.M[0] = 32'h010000EF;

    // Enter FETCH first (with reset asserted)
    wait_till_next_cfsm_state(FETCH);

    // Release reset
    reset = `FALSE;

    wait_till_next_cfsm_state(FETCH_WAIT);

    // -------- Single instruction: JAL x1, +16 --------

    // DECODE: verify opcode, rd and immediate
    wait_till_next_cfsm_state(DECODE);
    `assert_equal(uut.core.opcode, 7'b1101111)                    // JType (JAL)
    `assert_equal(uut.core.instruction_decode.rd,  5'd1)          // rd = x1
    `assert_equal(uut.core.instruction_decode.imm_ext, 32'sd16)   // imm = +16

    // UNCONDJUMP: link = pc_old + 4, PC updates by pc + imm
    wait_till_next_cfsm_state(UNCONDJUMP);
    `assert_equal(uut.core.alu.a, 32'd0)    // pc_old at address 0
    `assert_equal(uut.core.alu.b, 32'd4)
    `assert_equal(uut.core.alu.out, 32'd4)  // link value
    `assert_equal(uut.core.cfsm__pc_update, 1'b1)
    `assert_equal(uut.core.cfsm__pc_src, PC_SRC__JUMP)  // <-- enum literal, no hierarchy

    // ALUWB: write link back to rd (x1)
    wait_till_next_cfsm_state(ALUWB);

    // Back to FETCH: PC should be 16; x1 should be 4
    wait_till_next_cfsm_state(FETCH);
    wait_till_next_cfsm_state(FETCH_WAIT);
    `assert_equal(uut.core.RegFile.RFMem[1], 32'd4)  // rd = link = 4
    `assert_equal(uut.core.fetch.pc_cur, 32'd16)                                 // PC jumped to 16

    $finish;
  end

  `SETUP_VCD_DUMP(jal_only_tb)
/* verilator lint_off IMPORTSTAR */
/* verilator lint_off UNUSEDSIGNAL */
/* verilator lint_off INITIALDLY */

endmodule
