`include "src/types.svh"

module Mem_Stage (
    input wire RegWriteM,
    input logic [1:0] ResultSrcM,
    input wire MemWriteM,

);


endmodule