`include "src/types.svh"

module top ( input wire clk
           , input wire reset
           );

  wire     cfsm__pc_update;
  pc_src_t cfsm__pc_src;
  addr_t   pc_cur;
  addr_t   memory_address;
  data_t   data;
  instr_t  instruction;
  opcode_t opcode;
  imm_t    imm_ext;

  data_t __tmp_ResultData;

  data_t rd1;
  data_t rd2;

  data_t alu_input_a;
  data_t alu_input_b;

  addr_t pc_old;
  data_t Data; // TODO: this will need to be moved into fetch module

  wire alu__zero_flag;

  adr_src_t cfsm__adr_src;
  wire __tmp_IRWrite
     , __tmp_RegWrite
     , __tmp_MemWrite
     , __tmp_Branch;
  wire [1:0] __tmp_ALUSrcA
           , __tmp_ALUSrcB;
  wire [2:0] __tmp_ALUOp;
  wire [3:0] __tmp_ALUControl;
  wire [1:0] __tmp_ResultSrc;
  wire [3:0] __tmp_FSMState;
  data_t __tmp_ALUOut;

  ControlFSM control_fsm
    ( .opcode    ( opcode          )
    , .clk       ( clk             )
    , .reset     ( reset           )
    , .zero_flag ( alu__zero_flag  )
    , .AdrSrc    ( cfsm__adr_src   )
    , .IRWrite   ( __tmp_IRWrite   )
    , .RegWrite  ( __tmp_RegWrite  )
    , .PCUpdate  ( cfsm__pc_update )
    , .pc_src    ( cfsm__pc_src    )
    , .MemWrite  ( __tmp_MemWrite  )
    , .Branch    ( __tmp_Branch    )
    , .ALUSrcA   ( __tmp_ALUSrcA   )
    , .ALUSrcB   ( __tmp_ALUSrcB   )
    , .ALUOp     ( __tmp_ALUOp     )
    , .ResultSrc ( __tmp_ResultSrc )
    , .FSMState  ( __tmp_FSMState  )
    );

  fetch fetch
    ( .clk             ( clk             )
    , .reset           ( reset           )
    , .cfsm__pc_update ( cfsm__pc_update )
    , .cfsm__pc_src    ( cfsm__pc_src    )
    , .imm_ext         ( imm_ext         )

    // outputs
    , .pc_cur          ( pc_cur          )
    , .pc_old          ( pc_old          )
    );

  always @(*) begin
    case (cfsm__adr_src)
      ADR_SRC__PC:     memory_address = pc_cur;
      ADR_SRC__RESULT: memory_address = __tmp_ALUOut; // this will be the output of the result mux
    endcase
  end

  MA memory // instructions and data
    ( .A   ( memory_address )
    , .WD  ( 32'hxxxxxxxx   )
    , .WE  ( `FALSE         )
    , .CLK ( clk            )

    // outputs
    , .RD  ( data           )
    );

  Instruction_Decode instruction_decode
    ( .instr           ( data             )
    , .clk             ( clk              )
    , .reset           ( reset            )
    , .ResultData      ( __tmp_ResultData )
    , .opcode          ( opcode           )
    , .ALUControl      ( __tmp_ALUControl )
    , .baseAddr        ( rd1              )
    , .writeData       ( rd2              )
    , .imm_ext         ( imm_ext          )
    );

  ALU alu
    ( .a              ( rd1              )
    , .b              ( rd2              )
    , .alu_control    ( __tmp_ALUControl )
    , .out            ( __tmp_ALUOut     )
    , .zeroE          ( alu__zero_flag   )
    );

  always @(*) begin
    case (__tmp_ALUSrcA)
      ALU_SRC_A__PC:     alu_input_a = 32'd0;
      ALU_SRC_A__OLD_PC: alu_input_a = pc_old;
      ALU_SRC_A__RD1:    alu_input_a = rd1;
      default:           alu_input_a = 32'hxxxxxxxx;
    endcase
  end

  always @(*) begin
    case (__tmp_ALUSrcB)
      ALU_SRC_B__RD2:     alu_input_b = rd2;
      ALU_SRC_B__IMM_EXT: alu_input_b = imm_ext;
      ALU_SRC_B__4:       alu_input_b = 32'd4;
      default:            alu_input_b = 32'hxxxxxxxx;
    endcase
  end

  always @(*) begin
    case (__tmp_ResultSrc)
      2'b00: __tmp_ResultData = __tmp_ALUOut;
      2'b01: __tmp_ResultData = Data;
      2'b10: __tmp_ResultData = pc_old;
      default: __tmp_ResultData = 32'hxxxxxxxx;
    endcase
  end

endmodule
