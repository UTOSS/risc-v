`ifndef UTILS_VH
`define UTILS_VH

`define TRUE 1'b1
`define FALSE 1'b0

`endif
